module core #(
    parameter bw  = 4,       // bit-width of activations
    parameter col = 8,       // PE columns
    parameter row = 8,       // PE rows
    parameter psum_bw = 16,  // Partial sum bit-width 
    parameter ADDR_W = 11   // SRAM Address width
)(
    input                          clk,
    input                          reset,
    input [33:0]                   inst,           // 34-bit instruction packet from testbench
    input [bw*row-1:0]             D_xmem,         // Data written to x-mem by testbench
    output                         ofifo_valid,    // Write enable for FIFO output
    output [col*psum_bw-1:0]       sfp_out    // Output feature map
);

    wire acc;
    wire CEN_pmem;
    wire WEN_pmem;
    wire CEN_xmem;
    wire WEN_xmem;
    wire ofifo_rd;
    wire ififo_wr;
    wire ififo_rd;
    wire l0_rd;
    wire l0_wr;
    wire execute;
    wire load;

    wire [10:0] A_pmem;   // bits [30:20]
    wire [10:0] A_xmem;   // bits [17:7]

    assign acc       = inst[33];
    assign CEN_pmem  = inst[32];
    assign WEN_pmem  = inst[31];
    assign A_pmem    = inst[30:20];
    assign CEN_xmem  = inst[19];
    assign WEN_xmem  = inst[18];
    assign A_xmem    = inst[17:7];
    assign ofifo_rd  = inst[6];
    assign ififo_wr  = inst[5];
    assign ififo_rd  = inst[4];
    assign l0_rd     = inst[3];
    assign l0_wr     = inst[2];
    assign execute   = inst[1];
    assign load      = inst[0];

    wire [bw*row-1:0] Q_wt;

    sram #(
        .ADDR_W  (ADDR_W),
        .DATA_W (bw*row)   
    ) activation_sram (
        .CLK (clk),
        .CEN (CEN_xmem),
        .WEN (WEN_xmem),
        .A   (A_xmem),
        .D   (D_xmem),
        .Q   (Q_wt)
    );

endmodule
